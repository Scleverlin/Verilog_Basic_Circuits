// wait to start 

module TMUL_complex();

endmodule