module bf_tmul ();
input  





endmodule
