`include "/home/shi/verilog/FP_32/ADD_SUB/FP_32_add_or_sub.sv"
`include "/home/shi/verilog/FP_32/DIV/SRT_divider_FP32.sv"
`include "/home/shi/verilog/FP_32/MUL/FP32_mul.sv"
// RNE rounding mode
module FPU_32(op_code,a,b,result,clk,rst);




    

endmodule

