module post_processing(  //convert the final quotient to be IEEE-754
input logic [23:0] result,
input logic [4:0]shift_nums,
input logic right_shift,
input logic resultsign,
input logic [7:0] current_exponent,
output logic [31:0]quotient
);

logic [23:0] result_temp;
assign result_temp=(right_shift)?result>>shift_nums:result<<shift_nums;

logic [4:0] exponent_addend;
logic [23:0] result_shifted;

m_n_gen_2 mngen( result_temp,result_shifted,exponent_addend);
logic [7:0]exponent_final;

logic [7:0] addend_copmplement;

assign addend_copmplement=~exponent_addend+1;

assign exponent_final=current_exponent+addend_copmplement;

assign quotient={resultsign,exponent_final,result_shifted[22:0]};

endmodule


module m_n_gen_2 (
    input logic [23:0] data,
    output logic [23:0] outdata,
    output logic [4:0] shift
);
assign shift = (data[22] == 1) ? 0 :
               (data[21] == 1) ? 1 :
               (data[20] == 1) ? 2 :
               (data[19] == 1) ? 3 :
               (data[18] == 1) ? 4 :
               (data[17] == 1) ? 5 :
               (data[16] == 1) ? 6 :
               (data[15] == 1) ? 7 :
               (data[14] == 1) ? 8 :
               (data[13] == 1) ? 9 :
               (data[12] == 1) ? 10 :
               (data[11] == 1) ? 11 :
               (data[10] == 1) ? 12 :
               (data[9] == 1) ? 13 :
               (data[8] == 1) ? 14 :
               (data[7] == 1) ? 15 :
               (data[6] == 1) ? 16 :
               (data[5] == 1) ? 17 :
               (data[4] == 1) ? 18 :
               (data[3] == 1) ? 19 :
               (data[2] == 1) ? 20 :
               (data[1] == 1) ? 21 :
               (data[0] == 1) ? 22 : 0;

assign outdata = data << shift;
endmodule