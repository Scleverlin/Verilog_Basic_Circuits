// Prototype of shifterless Matrix-multiply design

module shifterLessFMA();

endmodule