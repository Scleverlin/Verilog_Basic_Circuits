// for easily changing the variable name