// wait to start 