module bf_tmul ();

endmodule
