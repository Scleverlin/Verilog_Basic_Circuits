// for easily changing the variable name


// multiplexer 0
extractor ex0  (sign_a,exp_a,RowB[0],RowC[0],sign_ab[0],exp_ab[0],sign_c[0],exp_c_minus_ab[0],mantissa_b[0],mantissa_c[0]);
extractor ex1  (sign_a,exp_a,RowB[1],RowC[1],sign_ab[1],exp_ab[1],sign_c[1],exp_c_minus_ab[1],mantissa_b[1],mantissa_c[1]);
extractor ex2  (sign_a,exp_a,RowB[2],RowC[2],sign_ab[2],exp_ab[2],sign_c[2],exp_c_minus_ab[2],mantissa_b[2],mantissa_c[2]);
extractor ex3  (sign_a,exp_a,RowB[3],RowC[3],sign_ab[3],exp_ab[3],sign_c[3],exp_c_minus_ab[3],mantissa_b[3],mantissa_c[3]);
extractor ex4  (sign_a,exp_a,RowB[4],RowC[4],sign_ab[4],exp_ab[4],sign_c[4],exp_c_minus_ab[4],mantissa_b[4],mantissa_c[4]);
extractor ex5  (sign_a,exp_a,RowB[5],RowC[5],sign_ab[5],exp_ab[5],sign_c[5],exp_c_minus_ab[5],mantissa_b[5],mantissa_c[5]);
extractor ex6  (sign_a,exp_a,RowB[6],RowC[6],sign_ab[6],exp_ab[6],sign_c[6],exp_c_minus_ab[6],mantissa_b[6],mantissa_c[6]);
extractor ex7  (sign_a,exp_a,RowB[7],RowC[7],sign_ab[7],exp_ab[7],sign_c[7],exp_c_minus_ab[7],mantissa_b[7],mantissa_c[7]);
extractor ex8  (sign_a,exp_a,RowB[8],RowC[8],sign_ab[8],exp_ab[8],sign_c[8],exp_c_minus_ab[8],mantissa_b[8],mantissa_c[8]);
extractor ex9  (sign_a,exp_a,RowB[9],RowC[9],sign_ab[9],exp_ab[9],sign_c[9],exp_c_minus_ab[9],mantissa_b[9],mantissa_c[9]);
extractor ex10 (sign_a,exp_a,RowB[10],RowC[10],sign_ab[10],exp_ab[10],sign_c[10],exp_c_minus_ab[10],mantissa_b[10],mantissa_c[10]);
extractor ex11 (sign_a,exp_a,RowB[11],RowC[11],sign_ab[11],exp_ab[11],sign_c[11],exp_c_minus_ab[11],mantissa_b[11],mantissa_c[11]);
extractor ex12 (sign_a,exp_a,RowB[12],RowC[12],sign_ab[12],exp_ab[12],sign_c[12],exp_c_minus_ab[12],mantissa_b[12],mantissa_c[12]);
extractor ex13 (sign_a,exp_a,RowB[13],RowC[13],sign_ab[13],exp_ab[13],sign_c[13],exp_c_minus_ab[13],mantissa_b[13],mantissa_c[13]);
extractor ex14 (sign_a,exp_a,RowB[14],RowC[14],sign_ab[14],exp_ab[14],sign_c[14],exp_c_minus_ab[14],mantissa_b[14],mantissa_c[14]);
extractor ex15 (sign_a,exp_a,RowB[15],RowC[15],sign_ab[15],exp_ab[15],sign_c[15],exp_c_minus_ab[15],mantissa_b[15],mantissa_c[15]);
