 module fast_lzc();

 endmodule;