module FMA_32();

endmodule
