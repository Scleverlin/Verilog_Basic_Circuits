// for easily changing the variable name


// multiplexer 0
